/*

*/



module #(parameter DATA_WIDTH = 8, SAMPLING =16)(
	input s_data_in,	
	input clk,reset,bclk,mode.
	output [DATA_WIDTH-1:0]p_data_out,
	output valid,
	output parity_error,stop_error);


endmodule
