`timescale 1ns/1ps

module tb_tx_control;

  // ------------------------------------------------------------
  // Parameters
  // ------------------------------------------------------------
  localparam CLK_FREQ   = 100_000_000; // 100 MHz
  localparam SAMPLING   = 16;
  localparam DATA_WIDTH = 8;

  // ------------------------------------------------------------
  // Testbench Signals
  // ------------------------------------------------------------
  reg clk;
  reg reset;
  reg ready;
  reg valid;
  reg [1:0] parity_select;
  reg [1:0] stop_select;
  reg [DATA_WIDTH-1:0] p_data_in;
  wire s_data_out;
  wire temp_busy;

  // ------------------------------------------------------------
  // DUT Instantiation
  // ------------------------------------------------------------
  uart_tx #(
    .DATA_WIDTH(DATA_WIDTH),
    .SAMPLING(SAMPLING)
  ) dut (
    .clk(clk),
    .reset(reset),
    .ready(ready),
    .valid(valid),
    .parity_select(parity_select),
    .stop_select(stop_select),
    .p_data_in(p_data_in),
    .s_data_out(s_data_out),
    .temp_busy(temp_busy)
  );

  // ------------------------------------------------------------
  // Clock Generation (100 MHz)
  // ------------------------------------------------------------
  initial begin
    clk = 0;
    forever #5 clk = ~clk; // 10 ns period -> 100 MHz
  end

  // ------------------------------------------------------------
  // Reset Task
  // ------------------------------------------------------------
  task apply_reset;
    begin
      reset = 1;
      valid = 0;
      ready = 0;
      @(posedge clk);
      @(posedge clk);
      reset = 0;
    end
  endtask

  // ------------------------------------------------------------
  // UART Transmission Stimulus
  // ------------------------------------------------------------
  task send_byte(
      input [DATA_WIDTH-1:0] data,
      input [1:0] parity_mode,
      input [1:0] stop_mode
  );
    begin
      @(posedge clk);
      parity_select = parity_mode;  // 00-none, 01-odd, 10-even
      stop_select   = stop_mode;    // 00-1 stop, 01-2 stops
      p_data_in     = data;
      valid         = 1;
      @(posedge clk);
      valid         = 0;
      $display("[%0t ns] Sending byte: 0x%0h (parity=%0b stop=%0b)", 
                $time, data, parity_mode, stop_mode);

      // Wait for transmission to complete
      wait (temp_busy == 1);
      wait (temp_busy == 0);
      $display("[%0t ns] Transmission complete.\n", $time);
    end
  endtask

  // ------------------------------------------------------------
  // Monitor serial output waveform
  // ------------------------------------------------------------
  initial begin
    $display("\n===== UART TX Testbench Start =====\n");
    apply_reset();

    // Test Case 1: No parity, 1 stop bit
    send_byte(8'hA5, 2'b00, 2'b00);

    // Test Case 2: Even parity, 1 stop bit
    send_byte(8'h3C, 2'b10, 2'b00);

    // Test Case 3: Odd parity, 2 stop bits
    send_byte(8'hF0, 2'b01, 2'b01);

    // Test Case 4: Random data
    send_byte(8'h55, 2'b00, 2'b00);

    $display("\n===== All UART TX Tests Completed =====\n");
    $finish;
  end


endmodule

