/*
Baud Generator 

*/

module baud_generator #(parameter SAMPLING = 16,CLK_FREQUENCY = 100000000, BAUD_RATA = 9600) (
	input clk,reset,
	output bclk);


endmodule
